module vmem(
    input               [9:0]       h_addr          ,
    input               [9:0]       v_addr          ,
    output              [23:0]      data_out        
);

assign data_out =   {8'd255, 8'd0, 8'd0};



endmodule
